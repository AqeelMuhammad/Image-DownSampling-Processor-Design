module instr_memory(
    input             clk, write_en,
    input      [15:0] addr, instr_in,
    output reg [15:0] instr_out
    );
    
    reg [15:0] ram [180:0];
    
    initial begin
	ram[0] = 8'd38;
	ram[1] = 16'd257;
	ram[2] = 8'd9;
	ram[3] = 8'd16;
	ram[4] = 8'd4;
	ram[5] = 8'd8;
	ram[6] = 8'd38;
	ram[7] = 8'd2;
	ram[8] = 8'd29;
	ram[9] = 8'd12;
	ram[10] = 8'd38;
	ram[11] = 8'd1;
	ram[12] = 8'd8;
	ram[13] = 8'd16;
	ram[14] = 8'd25;
	ram[15] = 8'd4;
	ram[16] = 8'd13;
	ram[17] = 8'd16;
	ram[18] = 8'd27;
	ram[19] = 8'd4;
	ram[20] = 8'd8;
	ram[21] = 8'd20;
	ram[22] = 8'd25;
	ram[23] = 8'd13;
	ram[24] = 8'd38;
	ram[25] = 16'd256;
	ram[26] = 8'd8;
	ram[27] = 8'd16;
	ram[28] = 8'd25;
	ram[29] = 8'd4;
	ram[30] = 8'd8;
	ram[31] = 8'd20;
	ram[32] = 8'd25;
	ram[33] = 8'd13;
	ram[34] = 8'd38;
	ram[35] = 16'd256;
	ram[36] = 8'd8;
	ram[37] = 8'd16;
	ram[38] = 8'd27;
	ram[39] = 8'd4;
	ram[40] = 8'd8;
	ram[41] = 8'd20;
	ram[42] = 8'd25;
	ram[43] = 8'd8;
	ram[44] = 8'd38;
	ram[45] = 8'd1;
	ram[46] = 8'd29;
	ram[47] = 8'd8;
	ram[48] = 8'd19;
	ram[49] = 8'd25;
	ram[50] = 8'd12;
	ram[51] = 8'd38;
	ram[52] = 16'd257;
	ram[53] = 8'd8;
	ram[54] = 8'd16;
	ram[55] = 8'd25;
	ram[56] = 8'd4;
	ram[57] = 8'd13;
	ram[58] = 8'd16;
	ram[59] = 8'd27;
	ram[60] = 8'd4;
	ram[61] = 8'd8;
	ram[62] = 8'd20;
	ram[63] = 8'd25;
	ram[64] = 8'd13;
	ram[65] = 8'd38;
	ram[66] = 8'd255;
	ram[67] = 8'd8;
	ram[68] = 8'd16;
	ram[69] = 8'd25;
	ram[70] = 8'd4;
	ram[71] = 8'd8;
	ram[72] = 8'd20;
	ram[73] = 8'd25;
	ram[74] = 8'd13;
	ram[75] = 8'd38;
	ram[76] = 8'd255;
	ram[77] = 8'd8;
	ram[78] = 8'd16;
	ram[79] = 8'd27;
	ram[80] = 8'd4;
	ram[81] = 8'd8;
	ram[82] = 8'd20;
	ram[83] = 8'd25;
	ram[84] = 8'd8;
	ram[85] = 8'd19;
	ram[86] = 8'd25;
	ram[87] = 8'd8;
	ram[88] = 8'd38;
	ram[89] = 8'd4;
	ram[90] = 8'd31;
	ram[91] = 8'd12;
	ram[92] = 8'd38;
	ram[93] = 16'd257;
	ram[94] = 8'd8;
	ram[95] = 8'd16;
	ram[96] = 8'd27;
	ram[97] = 8'd14;
	ram[98] = 8'd19;
	ram[99] = 8'd22;
	ram[100] = 8'd38;
	ram[101] = 16'd65278;
	ram[102] = 8'd8;
	ram[103] = 8'd16;
	ram[104] = 8'd27;
	ram[105] = 8'd41;
	ram[106] = 8'd127;
//	ram[106] = 8'd126;
	ram[107] = 8'd38;
	ram[108] = 8'd253;
	ram[109] = 8'd8;
	ram[110] = 8'd17;
	ram[111] = 8'd27;
	ram[112] = 8'd41;
	ram[113] = 8'd118;
	ram[114] = 8'd35;
	ram[115] = 8'd36;
	ram[116] = 8'd49;
	ram[117] = 8'd3;
	ram[118] = 8'd35;
	ram[119] = 8'd35;
	ram[120] = 8'd35;
	ram[121] = 8'd38;
	ram[122] = 8'd0;
	ram[123] = 8'd10;
	ram[124] = 8'd49;
	ram[125] = 8'd3;
	ram[126] = 8'd51;
	ram[127] = 8'd38;
	ram[128] = 8'd0;
	ram[129] = 8'd9;
	ram[130] = 8'd10;
	ram[131] = 8'd11;
	ram[132] = 8'd16;
	ram[133] = 8'd4;
	ram[134] = 8'd12;
	ram[135] = 8'd18;
	ram[136] = 8'd14;
	ram[137] = 8'd19;
	ram[138] = 8'd22;
	ram[139] = 8'd16;
	ram[140] = 8'd8;
	ram[141] = 8'd38;
	ram[142] = 16'd65278;
	ram[143] = 8'd27;
	ram[144] = 8'd41;
	ram[145] = 8'd172;
	ram[146] = 8'd17;
	ram[147] = 8'd8;
	ram[148] = 8'd38;
	ram[149] = 8'd254;
	ram[150] = 8'd27;
	ram[151] = 8'd41;
	ram[152] = 8'd160;
	ram[153] = 8'd36;
	ram[154] = 8'd36;
	ram[155] = 8'd35;
	ram[156] = 8'd35;
	ram[157] = 8'd37;
	ram[158] = 8'd49;
	ram[159] = 8'd132;
	ram[160] = 8'd38;
	ram[161] = 8'd0;
	ram[162] = 8'd10;
	ram[163] = 8'd38;
	ram[164] = 16'd258;
	ram[165] = 8'd8;
	ram[166] = 8'd16;
	ram[167] = 8'd25;
	ram[168] = 8'd9;
	ram[169] = 8'd37;
	ram[170] = 8'd49;
	ram[171] = 8'd132;
	ram[172] = 8'd51;
    end

    always @(posedge clk) begin
        if (write_en == 1)
            ram[addr] <= instr_in;
        else
            instr_out <= ram[addr];
        end
endmodule